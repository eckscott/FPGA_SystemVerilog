/***************************************************************************************
* 
* Filename: debounce_top.sv
*
* Author: Ethan Scott
* Description: connects the debounce module used to debounce a button
*              to the FPGA for the debouncing of one of the buttons on the
*              board
*
***************************************************************************************/
module debounce_top #(CLK_FREQUENCY=100_000_000, WAIT_TIME_US=5000,
                         REFRESH_RATE=200)(
    output logic[7:0] segment,      //7-seg display cathode seg outputs
    output logic[3:0] anode,        //7-seg display anode outputs
    input logic clk, btnd, btnc);   //clock, reset button, counter button

    logic sync_btnc;                 //synced button signals to global clock
    logic sync_btnc1;
    logic sync_reset1;
    logic sync_reset;             
    logic db_sig;                   //debounced signal
    logic pulse_out_db;             //output pulse generated by edge trigger
    logic pulse_out;
    logic f1_db, f2_db, f1, f2;     //intermediate flip flop vals used for edge trigger
    logic[7:0] counter_db;          //counts collective button pushes debounced
    logic[7:0] counter;             //counts collective button pushes not debounced

    logic[15:0] tot_count;          //total count that will be displayed with debounced
                                    //values being the lower 8 bits and undebounced being
                                    //the upper 8 bits
    localparam DP3_ON = 4'b0100;

    // Synce the button pushes to the global clock
    // sync 1
    always_ff @(posedge clk)
        sync_btnc1 <= btnc;
    // sync 2
    always_ff @(posedge clk)
        sync_btnc <= sync_btnc1;

    // sync 1
    always_ff @(posedge clk)
        sync_reset1 <= btnd;
    always_ff @(posedge clk)
        sync_reset <= sync_reset1;

    /******************************************* *
    * THE FOLLOWING IS FOR THE DEBOUNCED COUNTER *
    ******************************************* */
    // instantiating buttonDebouncer from the debounce module which connects everything
    // to the debouncer and debounces a button push
    debounce buttonDebouncer(.noisy(sync_btnc), .clk(clk), .rst(sync_reset),
                             .debounced(db_sig));

    // edge detector to verify one button push counts as 1 and doesn't increment 4ever
    // sync 1
    always_ff @(posedge clk)
        f1_db <= db_sig;
    // sync 2
    always_ff @(posedge clk)
        f2_db <= f1_db;
    // combination of 2 syncs
    assign pulse_out_db = (f1_db & ~f2_db);

    // Counter to count the button transitions
    always_ff @(posedge clk) begin
        if (btnd)
            counter_db <= 0;
        else if (pulse_out_db)
            counter_db <= counter_db + 1;
    end

    /********************************************* *
    * THE FOLLOWING IS FOR THE UNDEBOUNCED COUNTER *
    ********************************************* */
    // edge detector to verify one button push counts as 1 and doesn't increment 4ever
    always_ff @(posedge clk)
        f1 <= btnc;
    always_ff @(posedge clk)
        f2 <= f1;
    assign pulse_out = (f1 & ~f2);

    // Counter to count the button transitions
    always_ff @(posedge clk) begin
        if (btnd)
            counter <= 0;
        else if (pulse_out)
            counter <= counter + 1;
    end

    /********************************************* *
    *      CONNECT BOTH TO 7-SEGMENT DISPLAY       *
    ********************************************* */
    assign tot_count[7:0] = counter_db;
    assign tot_count[15:8] = counter;
    // instantiating sevenSegDisp as a module of a seven segment display to connect
    // these button pushes to be displayed on the seven segment display. Left 2 digits
    // showing debounced output and right 2 digits showing not debounced
    seven_segment4 sevenSegDisp(.segment(segment), .anode(anode), .data_in(tot_count),
                                .rst(btnd), .clk(clk), .dp_in(DP3_ON));

endmodule